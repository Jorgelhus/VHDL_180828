-- Projeto para dia 12 de Setembro:
-- Múltiplos de 5, exceto 0:
-- Saída 00
-- Valores: 5,10,15

-- Múltiplos de 3, exceto 0:
-- Pisca 1
-- Valores: 3,6,9,12

-- Múltiplos de 7, exceto 0:
-- Pisca 2
-- Valores: 7,14

-- Outros:
-- Aceso

-- Pisca 1 - 2x clock
-- Pisca 2 - 4x clock
-- 10 ciclos de clock